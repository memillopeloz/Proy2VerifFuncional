`ifndef SCOREBOARD_SV
`define SCOREBOARD_SV

class scoreboard;
	int dfifo[$]; // data fifo
	int afifo[$]; // address  fifo
	int bfifo[$]; // Burst Length fifo
endclass

`endif
