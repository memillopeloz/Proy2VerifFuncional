class transaction;
	logic bl;
	logic address;
	logic value;
endclass
