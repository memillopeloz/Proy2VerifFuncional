`ifndef TEST_1_SV
`define TEST_1_SV

program test_1(sdrc_if sdrc_intf);
	initial begin
		$display("-------------------------------------- ");
		$display(" Case-1: Single Write/Read Case        ");
		$display("-------------------------------------- ");
	end
endprogram

`endif