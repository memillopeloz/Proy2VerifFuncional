`ifndef TRANSACTION_SV
`define TRANSACTION_SV

class transaction;
	logic bl;
	logic [32:0] address;
	logic value;
endclass

`endif