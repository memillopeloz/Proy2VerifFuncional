`ifndef TRANSACTION_SV
`define TRANSACTION_SV

class transaction;
	logic [32:0] address;
	logic bl;
	logic value;
endclass

`endif